//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-6
//Part Number: GW5A-LV25MG121NES
//Device: GW5A-25
//Device Version: A
//Created Time: Sat Dec 09 13:40:27 2023

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire [23:0] prom_inst_1_dout_w;
wire [23:0] prom_inst_2_dout_w;
wire [23:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h68E527C2775F5FB90FEB31DBB71E3F1F3E3E3FFD9A799A9A9A9A9A9A977495D7;
defparam prom_inst_0.INIT_RAM_01 = 256'h9A9A9A9A9A999A9A9A9A9A9A9A9A9A9A9A9ABABABABABABBBBBBBABBBB080BEB;
defparam prom_inst_0.INIT_RAM_02 = 256'h870405C436FE738586C725CAC7703E3F3F1D9B999A9A9A9A9A9A9A997595B6B6;
defparam prom_inst_0.INIT_RAM_03 = 256'h9A9A9A9A9A9A9A9BBABA9A9A9A9B9A9ABABBBA9A9A9A9ABBBBBABABBBB080BEB;
defparam prom_inst_0.INIT_RAM_04 = 256'h8948E58FDBB8ED43478A4D480888343FDC9A9A9A9A9A9A9A9A9AB97595B6B6B6;
defparam prom_inst_0.INIT_RAM_05 = 256'h9A9A9A9A9A9BBBBA97779777B9BBBBBBBBBBBA9A9A9A9ABABBBBBABB9A07EA0C;
defparam prom_inst_0.INIT_RAM_06 = 256'h2626A391B774F88C8407086BC7C755BC7A9A9A9A9A9A9A9A9BBB9794B5B6B6B6;
defparam prom_inst_0.INIT_RAM_07 = 256'h9A9A9A9A9ABABA987474747476BBBBBBBBBA9A9A9A9A9A9ABABABABB9A07EA2D;
defparam prom_inst_0.INIT_RAM_08 = 256'h8946A26D96D71868C62806EB48E931BB9C9A9A9A9A9A9A9ABA9875B6B6B6B6B6;
defparam prom_inst_0.INIT_RAM_09 = 256'h9A9A9A9ABA9BB9757494747475B9BBBB9A9A9A9B999B9A999A9BBADBBB08EAEB;
defparam prom_inst_0.INIT_RAM_0A = 256'h896783AC18B6F00724C8E7484CE94410BB9B9A9A9A9A9ABA9795B6B6B6B6B696;
defparam prom_inst_0.INIT_RAM_0B = 256'h9A9A9ABA9A9B9875947575757475B9BA9A9BBB9B999B9ABB9A9A9BBCBB08EB88;
defparam prom_inst_0.INIT_RAM_0C = 256'h6867066A314A694881A528A6C56345EF9799BA9A9B9B9A9775B5B6B6B6B6B695;
defparam prom_inst_0.INIT_RAM_0D = 256'h9A9ABABA9A997674747575757575757698BA9B9BBBBC9A56BC9C9ABABB08EBA9;
defparam prom_inst_0.INIT_RAM_0E = 256'h6889A9486ACB6769ABE2A3A5E4AE9796757598BA9B9A9875B5D6B6B6B6B69696;
defparam prom_inst_0.INIT_RAM_0F = 256'h9ABABA9A9A96747475757575757574747597BB577654CDA7AE7ABABABB080CEC;
defparam prom_inst_0.INIT_RAM_10 = 256'h468988EA0CE548B7B8ADA20105757594947595989A987596B6B6B7B6B6B6B696;
defparam prom_inst_0.INIT_RAM_11 = 256'hBABA9A9A997574747575757575759494749495EB0B4847E905CA99BD9A080CEC;
defparam prom_inst_0.INIT_RAM_12 = 256'h26680547271195B67696528B1095947474757575969596B6B6B6B6B6B6B5B6B5;
defparam prom_inst_0.INIT_RAM_13 = 256'h9A9A9ABA7674747575757575757595947573A8C987E6892B684579BB9B07EBEB;
defparam prom_inst_0.INIT_RAM_14 = 256'h8805C5C551F7D69575769594B6957575759595757495B6B6B6B6B6B6B5B6B695;
defparam prom_inst_0.INIT_RAM_15 = 256'h9A9A99977574757575757575757575947595A9064D480BAA6434BBBB9A07CA0D;
defparam prom_inst_0.INIT_RAM_16 = 256'hA946C4AD17D6B595757595B6D7B7B5757595759596B6B6B6B6B6B6B5B6B6B695;
defparam prom_inst_0.INIT_RAM_17 = 256'h9A9876757475757575757575757574749695EBE7482889E62457DBBA76060C2D;
defparam prom_inst_0.INIT_RAM_18 = 256'h6788A3ADF8B69574947495B6B6B6B69574959596B6B6B6B6B6B6B6B6B6B69575;
defparam prom_inst_0.INIT_RAM_19 = 256'h96757475757575757575757575757474968C04E74264E785A22999B79506EBEC;
defparam prom_inst_0.INIT_RAM_1A = 256'hA947A2ADF8B69574747495B6B6B69575749596B6D6B6B6D6B6B6B6B6B6B69574;
defparam prom_inst_0.INIT_RAM_1B = 256'h94947475757575757574747575959595956AC001C62AE801A28A4AAC3106EB0C;
defparam prom_inst_0.INIT_RAM_1C = 256'hEB27C4ADF8B675757595B6B6B6B6757475759595B6B6D6B695959595B5957475;
defparam prom_inst_0.INIT_RAM_1D = 256'h75757575747575757575959575959596B5B5AC4685E622E68C48A8AB29890B2C;
defparam prom_inst_0.INIT_RAM_1E = 256'h8905068CD895747495B6B6B6B6B675747495957475959595B6B6B69574757575;
defparam prom_inst_0.INIT_RAM_1F = 256'h757575757575757575747575747574759595D912E2E0E3F1D7CDC5482D2C2CEC;
defparam prom_inst_0.INIT_RAM_20 = 256'h4626C48CD7957495B6B6B6B6B6B69595959575757575749595B6B6B695757575;
defparam prom_inst_0.INIT_RAM_21 = 256'h75757575757575757575757575757575757596936AAC32B47595528C27890CEB;
defparam prom_inst_0.INIT_RAM_22 = 256'h4647C48DF89595B6B6B6B6B6B6B69595B67475957495B596959595B6B6957575;
defparam prom_inst_0.INIT_RAM_23 = 256'h75757575757575757575757574759574747495959595B674767595B6ADA50CE9;
defparam prom_inst_0.INIT_RAM_24 = 256'hAA26C4ADD996B6B6B6B6B6B6B6B6957595957575757595B6B6B6B69595957574;
defparam prom_inst_0.INIT_RAM_25 = 256'h757575757575757574959574957475757474757595957475957574959527EA0D;
defparam prom_inst_0.INIT_RAM_26 = 256'h8989E48BD7B6D6B6B6B6B6B6B6B6B575959595757575749495B6B6B6B6B69595;
defparam prom_inst_0.INIT_RAM_27 = 256'h7575757575757575759595759595747575757575757575757475759595E6A92D;
defparam prom_inst_0.INIT_RAM_28 = 256'hA96905E531D6D6B6B6B6B6B6B6B695757595959595959595949495B6B6B6D6B6;
defparam prom_inst_0.INIT_RAM_29 = 256'h75757575757575757574757475B695949575747575757575757575B6AD06AA2C;
defparam prom_inst_0.INIT_RAM_2A = 256'hCA264726A5B5D7B6B6B6B6B6B6B69574757475959595959595957495959595B6;
defparam prom_inst_0.INIT_RAM_2B = 256'h7575757575757575757575759595B6B595747475757475757575957327A80DEC;
defparam prom_inst_0.INIT_RAM_2C = 256'hCA480547C4ACD7D7B6B5D5D6B595957474757574747574757495B69474747595;
defparam prom_inst_0.INIT_RAM_2D = 256'h7574749575759594759475959475B5D6B5747575949594749575D8AE476ECBAA;
defparam prom_inst_0.INIT_RAM_2E = 256'hA968058A05A5D6D7F8B796957576949474947594737595B5B59494B595947574;
defparam prom_inst_0.INIT_RAM_2F = 256'h74949475747574947574757474747496D6B575747475759594736B4A0C2C0BEB;
defparam prom_inst_0.INIT_RAM_30 = 256'h88680648680605E731F796D6B69695967694977696B6B7D6D8B5959797B69575;
defparam prom_inst_0.INIT_RAM_31 = 256'hD6D7D9D8D6B7969696969595989596D7D7B7D67596B6B7EF0847EB0CEBEB2D2D;
defparam prom_inst_0.INIT_RAM_32 = 256'hCAC4A447682727A36352FB7497EF52147673AF7511CE76F733F933CD13D83196;
defparam prom_inst_0.INIT_RAM_33 = 256'hF975F111F875953233545476B05412CD751932F854CE8D280D474867058AED68;
defparam prom_inst_0.INIT_RAM_34 = 256'hA7E6268782A7A56447E98E0AAC27E9CBAAAA27CAE826CB8CE98DCA24EA6BE9AB;
defparam prom_inst_0.INIT_RAM_35 = 256'h6DCA26088CCB09E9EAEAACAA27CCE825CB8CE98CCB46C6C3C8E3068546A38847;
defparam prom_inst_0.INIT_RAM_36 = 256'hA96CCD0AC96B874BCD4B674AE98B2A2BE8EA4BA98BADEBA84B872BAC4C886CC9;
defparam prom_inst_0.INIT_RAM_37 = 256'h670ACD8D872A094C4B0AEAE84B684BADEBA86C880AAD8C892A2A8C4B4CEAEA2C;
defparam prom_inst_0.INIT_RAM_38 = 256'h056DEB464B6CADC8660A670B6D47EAC9882BE5478CCA474B6C8DC826470A6C8C;
defparam prom_inst_0.INIT_RAM_39 = 256'hCDEA270B87CA6D67C9EA874C05066C0C472A4CAEC9260A67CA6C47E9C8872CC5;
defparam prom_inst_0.INIT_RAM_3A = 256'h84AAE644C567CA6464E645C60765E5A665C64584EBC624C688CA852545A626EA;
defparam prom_inst_0.INIT_RAM_3B = 256'hEAC664C664A60785A5C665C76564AA2744A548EBC544E645A62845C5A544C665;
defparam prom_inst_0.INIT_RAM_3C = 256'h678545894665856768668966456865886846A966A587894685A56889894765C5;
defparam prom_inst_0.INIT_RAM_3D = 256'h8566A845A96744884566884689678566896665A5678946A967458844678846A9;
defparam prom_inst_0.INIT_RAM_3E = 256'h8946A9AA8A6847AAA989A9A988896889A989AA894689AAA96847AAA9A9898947;
defparam prom_inst_0.INIT_RAM_3F = 256'h47A9A989AAA988A988A8A9A9AAA96788A9A968468AAA89A9A989A98889A9A9A9;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[23:0],dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 8;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h3D28392042575B3A26152E463A53534F53534F42363636363636363A322A2A2A;
defparam prom_inst_1.INIT_RAM_01 = 256'h36363636363A3A36363636363636363636363636363636363636363636255A55;
defparam prom_inst_1.INIT_RAM_02 = 256'h413131182E4232050A12021909265753534B3A3636363636363636362A2A2A2A;
defparam prom_inst_1.INIT_RAM_03 = 256'h36363636363636363636363636363636363A3636363636363636363636215A55;
defparam prom_inst_1.INIT_RAM_04 = 256'h453D2C2D362A19050E0E0F0E0F0232533E363636363636363636362A262A2A2A;
defparam prom_inst_1.INIT_RAM_05 = 256'h36363636363636362E2E2E2E363636363A363636363636363A3636363621555A;
defparam prom_inst_1.INIT_RAM_06 = 256'h3535242932262E15050E0E0E0A092E3E363636363636363636362E262A2A2A2A;
defparam prom_inst_1.INIT_RAM_07 = 256'h363636363636362E2A26262A2E3A36363636363636363636363636363621555E;
defparam prom_inst_1.INIT_RAM_08 = 256'h453524252E2A27150D12060E0E0D263A363636363636363A362E262A2A2A2A2E;
defparam prom_inst_1.INIT_RAM_09 = 256'h363636363636362A2626262A2A363A363636363A3A3A36363A3A363636255555;
defparam prom_inst_1.INIT_RAM_0A = 256'h493D24212B262531150D0D0E130E09223A3A3A363636363A2E2A2A2A2A2A2E2A;
defparam prom_inst_1.INIT_RAM_0B = 256'h36363636363A322A26262A2A262A3636363A3636363636363636363636255545;
defparam prom_inst_1.INIT_RAM_0C = 256'h454135212221414910010E0D05090D1D32363A3A3A3A362E2A2A2A2A2A2A2A26;
defparam prom_inst_1.INIT_RAM_0D = 256'h3636363636362E2A2A262A262A2A2A2E3236363A363A3A363A32363A36215949;
defparam prom_inst_1.INIT_RAM_0E = 256'h4545413941554929190405090421322A2A2E32363A3A2E262A2E2A2A2A2A2A2A;
defparam prom_inst_1.INIT_RAM_0F = 256'h36363A3A362E2A2A2A2A2A2A2A2A2A2A2A2E3E362E2619151D363A3636255E55;
defparam prom_inst_1.INIT_RAM_10 = 256'h39494951563021222A1D0805052E2A2626262A323A32262A2A2A2A2A2A2A2A2A;
defparam prom_inst_1.INIT_RAM_11 = 256'h3636363A362A2A2A2A2A2A2A2A2A262A2A2A32150E0E0E060619363636255E55;
defparam prom_inst_1.INIT_RAM_12 = 256'h3939353D25262A262A2A2A15222A262A2A2A262A2E2A2A2A2A2A2A2E2A2A2A26;
defparam prom_inst_1.INIT_RAM_13 = 256'h363636362E262A2A2A2A2A2A2A26262A2A2A0D0A0611120F0E0D3A3636255955;
defparam prom_inst_1.INIT_RAM_14 = 256'h41352C182E322A262A2A2A2E2E26262A2A262A2A262A2E2A2A2A2A2A2A2A2A26;
defparam prom_inst_1.INIT_RAM_15 = 256'h3A36362E26262A2A2A2A2A2A2A2A2A26262A0D0A1B0A0F12012A3E363221555A;
defparam prom_inst_1.INIT_RAM_16 = 256'h453D28252B2A2A262A2A262A2A2A2A2A2A2626262A2A2A2A2A2A2A2A2A2A2A2A;
defparam prom_inst_1.INIT_RAM_17 = 256'h36322A26262A2A2A2A2A2A2A2A2A2A26262E1909120E0E09052E3A362A215A5E;
defparam prom_inst_1.INIT_RAM_18 = 256'h414524212A2E2A26262A2A2A2A2A2A262626262A2A2A2A2A2A2A2A2A2A2A2A2A;
defparam prom_inst_1.INIT_RAM_19 = 256'h2A2A262A2A2A2A2A2A2A2A2A2A2A2A2A2E19050D0505090910213A32261D5559;
defparam prom_inst_1.INIT_RAM_1A = 256'h4D3D20212E2E2A2A2A2A2A2A2A2A2A2A262A2A2A2A2A2A2A2A2A2A2A2A2A2626;
defparam prom_inst_1.INIT_RAM_1B = 256'h26262A2A2A2A2A2A2A26262A2A2A26262E1500050912090524452D21221D555A;
defparam prom_inst_1.INIT_RAM_1C = 256'h553928252A2A2A2A2A262A2A2A2A2A262A2A2A262A2A2A2A262A2A2A2A2A262A;
defparam prom_inst_1.INIT_RAM_1D = 256'h2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A262A321D0D050D01102131554D3545565A;
defparam prom_inst_1.INIT_RAM_1E = 256'h493131252A2A26262A2A2A2A2A2A2626262A2A2A2A2A2A2A2A2E2E2A262A2A2A;
defparam prom_inst_1.INIT_RAM_1F = 256'h2A2A2A2A2A2A2A2A2A262A2A262A2A2A2A2A3226040404252E2124415E5A5A59;
defparam prom_inst_1.INIT_RAM_20 = 256'h3D3528252A2A26262A2A2A2A2A2A2A262A2A2A2A2A2626262A2A2E2E2A2A2A2A;
defparam prom_inst_1.INIT_RAM_21 = 256'h2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A26262A151D26262A2E1E2139495E55;
defparam prom_inst_1.INIT_RAM_22 = 256'h393928252E2A2A2A2A2A2A2A2A2A26262A26262626262A2A2A2A2A2A2A262626;
defparam prom_inst_1.INIT_RAM_23 = 256'h2A2A2A2A2A2A2A2A2A2A2A2A2626262A2A2A262A2A2A2A2A262A2E2A21205A51;
defparam prom_inst_1.INIT_RAM_24 = 256'h45352C212A2A2A2E2A2A2A2A2A2A262A2A2A262A26262A2A2A2A2A2A2A2A2626;
defparam prom_inst_1.INIT_RAM_25 = 256'h2A2A2A2A2A2A2A2A262A2A262A262A2A2A2626262A26262A262A2A262219555E;
defparam prom_inst_1.INIT_RAM_26 = 256'h45452C212E26262E2A2A2A2A2A2A2A2A2A2A2A2A2A2A26262A2A2E2E2E2A2A26;
defparam prom_inst_1.INIT_RAM_27 = 256'h2A2A2A2A2A2A2A2A2A2A2A262A2A262A2A2A2A2A2A2A2A262A2A2A26261C515A;
defparam prom_inst_1.INIT_RAM_28 = 256'h4941311C2A2E262A2A2A2A2A2A2A262A2A2A2A2A2A2A2A2626262A2A2A2A2A2A;
defparam prom_inst_1.INIT_RAM_29 = 256'h2A2A2A2A2A2A2A2A2A262626262E2A262A2A2A2A2A2A2A2A2A2A262A1D31515A;
defparam prom_inst_1.INIT_RAM_2A = 256'h4D353935102A2A2A2A2A2A2A2A2A26262A26262A2A2A2A2A2A2626262A2A2A2A;
defparam prom_inst_1.INIT_RAM_2B = 256'h2A2A2A2A2A262A2A2A2626262A2A2A2A262A2A2A2A2A2A2A2A262A2A2D495A59;
defparam prom_inst_1.INIT_RAM_2C = 256'h4D3D353D20252E2E2E2A2A2A2A2A262E2A2A262A2A2A2A2A2A2A2A26262A2A26;
defparam prom_inst_1.INIT_RAM_2D = 256'h2A262626262A2626262626262626262A2A2A262A2626262A2A2E261D41665551;
defparam prom_inst_1.INIT_RAM_2E = 256'h453D2D45351C262A262E2E262A2A26262A2626262A2A262A262A2A2A2A262A2A;
defparam prom_inst_1.INIT_RAM_2F = 256'h2A2A2A2A2A2A26262A2A2A26262E2A2E2A2A2A2A262A2E261E2A19355A5A5651;
defparam prom_inst_1.INIT_RAM_30 = 256'h493D2D4149351D242A2A2A2A2A2E2E222A2A2A2A2A2A2A2A2E2A2A2A2A262A2E;
defparam prom_inst_1.INIT_RAM_31 = 256'h262A2E2E26262A2A2A262A262E26262A262E2A2A2A2626252D2D555E5559565E;
defparam prom_inst_1.INIT_RAM_32 = 256'h512C243541393928181E2E2A2E1D262A2A2625261E1D2A2E262E2215262A2226;
defparam prom_inst_1.INIT_RAM_33 = 256'h322A21222E2A2E222A262A2E1D2626192A2B2A262A1D15455E414939314D5D45;
defparam prom_inst_1.INIT_RAM_34 = 256'h1D110621180D240D060D1D1215060D15151106150D02151D0D19110609190D11;
defparam prom_inst_1.INIT_RAM_35 = 256'h1D11020E1915120D111111150A150D0215190D191102091C210C060909142D06;
defparam prom_inst_1.INIT_RAM_36 = 256'h0A0B0F0F060B0A0F0F130A0B0A130F0B06120F0E0B130A0A0B06131313060B0E;
defparam prom_inst_1.INIT_RAM_37 = 256'h0A0B0B130A0B0B130B0F0E0613120B130E060F0A0B0F130E070F0F0F0B060A0F;
defparam prom_inst_1.INIT_RAM_38 = 256'h0A0F12060B13130A060B060F0F060E0E0A0B01060F12020B13130E02020B1313;
defparam prom_inst_1.INIT_RAM_39 = 256'h0B120613060E13060A0E060F06060F0F0A0B13130A0A0B0A0E130A0A06060F05;
defparam prom_inst_1.INIT_RAM_3A = 256'h0D0E111D11060E19190D1D150E1505151D111D0D0A112115060A15211D15060A;
defparam prom_inst_1.INIT_RAM_3B = 256'h06151D1519150A1509111D15190D0E0A1D150A0A1121111D190A190915211119;
defparam prom_inst_1.INIT_RAM_3C = 256'h3111294D3119153D49314935293D21394135492D0D314D351911394D493D1D0D;
defparam prom_inst_1.INIT_RAM_3D = 256'h1131453141352539293545314535152949311D113549354535253D293D453145;
defparam prom_inst_1.INIT_RAM_3E = 256'h4D39494D5145394D514D5149494D4D51514D4D49354D5149413D4D4D51514931;
defparam prom_inst_1.INIT_RAM_3F = 256'h3549514D4D4D494D494D4D495149354D55494535514D4D514D4D4D494D4D4951;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[23:0],dout[23:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 8;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h5F7F7F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F;
defparam prom_inst_2.INIT_RAM_01 = 256'h9EBFBFBF7E5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5E5F5F;
defparam prom_inst_2.INIT_RAM_02 = 256'h5F7E5F5F7F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F;
defparam prom_inst_2.INIT_RAM_03 = 256'hBEBFBFBFBFBF7E5E5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F7F5F5F7F5E;
defparam prom_inst_2.INIT_RAM_04 = 256'h7F5F5F7E7E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_2.INIT_RAM_05 = 256'hBFBFBFBFBFDFBE9E9F9F7E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7E7E7F7F7F;
defparam prom_inst_2.INIT_RAM_06 = 256'h7EADB07F5F7F9F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_2.INIT_RAM_07 = 256'hBFBF9EBFBFBFBFDFDFBE9F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F5D8BF4;
defparam prom_inst_2.INIT_RAM_08 = 256'h634505F3BF7F3B3B7F9F7F7E7E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_2.INIT_RAM_09 = 256'hDFBFBFBFBFBFBFDFDEDEDF9F7F7F7E7E7F7F7F7F7F7F7F7F7F7F3B7E7E6805C6;
defparam prom_inst_2.INIT_RAM_0A = 256'hA60627AD37F12384D0399F7F7E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_2.INIT_RAM_0B = 256'hDFDFDFDFDEDEBEBEBEBFBFBF9F9F9EBFDFBF9E7F7F7F7F7FBF3785CE6EA5886A;
defparam prom_inst_2.INIT_RAM_0C = 256'hE7E66A27C5624747A26615BF7F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F;
defparam prom_inst_2.INIT_RAM_0D = 256'hDFDFDFBCBBBBBCBD9D9F9F7F7F7EDEDFDFDFBE9E9F7F7FBF38C448A4C56868E7;
defparam prom_inst_2.INIT_RAM_0E = 256'hA9EACACA680669496A2645399F9E9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F;
defparam prom_inst_2.INIT_RAM_0F = 256'hDFFFBC9ABADABBBB9C9D9EBFDFDFDFDEDFDEDFDF9E9EBF5A25486B460A0D8AE7;
defparam prom_inst_2.INIT_RAM_10 = 256'hAA0A2BAA690BEB27276843F3BF9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F;
defparam prom_inst_2.INIT_RAM_11 = 256'hFEBC9ABBBBBBBBBBBABA9ADDFFFFDFDFFFDFDFFFDFDFFFF2824767CBEB87EA2C;
defparam prom_inst_2.INIT_RAM_12 = 256'hCAC96BCA4889AB0785834759BF9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F;
defparam prom_inst_2.INIT_RAM_13 = 256'hBB9ABABBBBBBBBBA9A9A9A9ADDFEDFDFDFFFFFFEFF1F1584ABC6274DAAA9A8EB;
defparam prom_inst_2.INIT_RAM_14 = 256'h6A4D2B69CBAACAE6E6628FDFBEDFBF9F9F9FBFBFBFBFBFBFBFBFBFBFBFBFBFBF;
defparam prom_inst_2.INIT_RAM_15 = 256'h9ABABABBBBBA9A9A9A9A9A9A9ADDFFFFDFDFDFDF1F1403A48B690669690CEBE7;
defparam prom_inst_2.INIT_RAM_16 = 256'h484788698A2CEB8A27A304573FFFFFBEBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBF;
defparam prom_inst_2.INIT_RAM_17 = 256'hBBBBBABBBB9A9A9A9A9A9A9A9A9ADDFFDEBFDFFF9D4A25E68469EB8927C5698A;
defparam prom_inst_2.INIT_RAM_18 = 256'hA967A92C692748E7A50764D0BC1FFFFFDFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBF;
defparam prom_inst_2.INIT_RAM_19 = 256'hBBBBBBBBBB9A9A9A9A9A9A9A9A9A9A9CBFBFBF14E4238A49C4262CEB89E6CA2C;
defparam prom_inst_2.INIT_RAM_1A = 256'h0C4C88AA682727E608C6A64203531F1FFFDFDFDFDFBFBFBFBFBFBFBFBFBFBFBF;
defparam prom_inst_2.INIT_RAM_1B = 256'hBBBBBBBBBA9A9A9A9A9A9A9A9A9A9A7BBDFF5AC2C384A5480B0B680CEA488AEB;
defparam prom_inst_2.INIT_RAM_1C = 256'h276869E7078AEB0B89268B07206A1F1F1FFEFF1FFFDFBFBFBFBFBFBFBFBFBFDF;
defparam prom_inst_2.INIT_RAM_1D = 256'hBBBBBBBABA9A9A9A9A9A9A9A9A9A9A9A9ABBBED24464238348EA0668CAAA6928;
defparam prom_inst_2.INIT_RAM_1E = 256'h07A489EBCA48EBA9280BEAA48CBC1F1FFF1F1F1FFFFFDEDFDFDFDFDFDFDFDFDF;
defparam prom_inst_2.INIT_RAM_1F = 256'hBBBBBBBABA9A9A9A9A9A9A9A9A9A9A9A9A9ABCFF8FA6E7648427A9EAEBCA88A9;
defparam prom_inst_2.INIT_RAM_20 = 256'hEB0727A92C0B4808E728A6E2341FFFFFFFFFFFFFFFFFFFDFDFDFDFDFDFDFDFDF;
defparam prom_inst_2.INIT_RAM_21 = 256'hBBBBBBBA9A9A9A9A9A9A9A9A9A9A9A9A9A9ABC34E2E7E744438427EBA947A90B;
defparam prom_inst_2.INIT_RAM_22 = 256'hEBA92CEB68A98A49C6848686E3F4FFDFDFDFDFDFDFFFDFDFDFDFDFDFDFDFDFFF;
defparam prom_inst_2.INIT_RAM_23 = 256'hBBBBBBBA9A9A9A9A9A9A9A9A9A9A9A9A9A9ABB7A6B21A6A6C6E8A58428CBCBA9;
defparam prom_inst_2.INIT_RAM_24 = 256'hA506CC8AA5A4C78584E7C684236DFFDFDFDFDFDFDFDFDFDEDEDFDFDFDFDFFF1F;
defparam prom_inst_2.INIT_RAM_25 = 256'hBBBBBBBA9A9A9A9A9A9A9A9A9A9A9A9A9A9ABB570843E728E7084A2806484D69;
defparam prom_inst_2.INIT_RAM_26 = 256'hA5A5E7E707286485286A2640069BFFFFDFDFDFDFDFDFDFDFDFDFDFDFFFFF1F1F;
defparam prom_inst_2.INIT_RAM_27 = 256'hBBBBBB9A9A9A9A9A9A9A9A9A9A9A9A9A9A9ABD11A045848364A5E749AA6948C5;
defparam prom_inst_2.INIT_RAM_28 = 256'h280807288B28A5A528084464014A1FFFFFFFFFFFFFFFFFDFFFDFFF1F1F1F1E1E;
defparam prom_inst_2.INIT_RAM_29 = 256'hBBBABA9A9A9A9A9A9A9A9A9A9A9A9A9A9A9ABB5627238429A5C60808E6088A48;
defparam prom_inst_2.INIT_RAM_2A = 256'h288B49C5C643A528A584A420E4571FFFFFFFFFFFFFFFFFFFFFFF1F1F1F1F1F1F;
defparam prom_inst_2.INIT_RAM_2B = 256'hBABA9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A99DDB0C06508A50828C6C643C608;
defparam prom_inst_2.INIT_RAM_2C = 256'hC6E7C5E764A56A49A5C4C5E4561FFFFFFFFFFFFFFFFFFFFF1F3F1E1E1F1F1F1F;
defparam prom_inst_2.INIT_RAM_2D = 256'hBBBBBABA9A9A9A9A9A9A9A9A9A9A9A9A9A9A9B9C780622854384A784E7082284;
defparam prom_inst_2.INIT_RAM_2E = 256'hC68464C7C6A5E7864400E02AFE1FFFFFFFFFFFFFFF1F1F3E3F3F1E1E3F3F3F3F;
defparam prom_inst_2.INIT_RAM_2F = 256'hBBBABABA9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9BBCAEC1E163E6C642C6084264;
defparam prom_inst_2.INIT_RAM_30 = 256'hE7432364A54342E4456E6E991FFF1F1F1F1F1F1F1F1F1F1F1F1F1E1E1F1F1F3F;
defparam prom_inst_2.INIT_RAM_31 = 256'hBA9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9BBBAF2722C700A20301C385;
defparam prom_inst_2.INIT_RAM_32 = 256'h65E223C6C602E260261E5F1F1F1F1F1F1F1F1F1F1F1F1F1E1E1F1F1E1E1E1E1E;
defparam prom_inst_2.INIT_RAM_33 = 256'h9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9B9BDC9B2BA214584AA1C524;
defparam prom_inst_2.INIT_RAM_34 = 256'hC3A30364E08B1406763F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F;
defparam prom_inst_2.INIT_RAM_35 = 256'h9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A99999ABC7A37FE7FFC0947E4;
defparam prom_inst_2.INIT_RAM_36 = 256'hE506C3074DFD3F1E3F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F;
defparam prom_inst_2.INIT_RAM_37 = 256'h9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A99BBBD9ADC3F4A8726;
defparam prom_inst_2.INIT_RAM_38 = 256'h260682F29F3F1F3F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F3F3F3F3E;
defparam prom_inst_2.INIT_RAM_39 = 256'h9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9ABC29CAAA;
defparam prom_inst_2.INIT_RAM_3A = 256'h674782F25F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F3F1F1F1F1FFDFDFC98;
defparam prom_inst_2.INIT_RAM_3B = 256'h9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9ABB9A080CAA;
defparam prom_inst_2.INIT_RAM_3C = 256'h680505E8995F3F1F1F3F1F1F1F1F1F1F1F1F1F1F3F3F3FFDBB9A9A9A7A9A7674;
defparam prom_inst_2.INIT_RAM_3D = 256'h9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9ABBBB08EBEC;
defparam prom_inst_2.INIT_RAM_3E = 256'h69E405C4775F1F5F3FBC5F3F3F3F1F1F1F1F3F3F1EDD9B9A9A9A9A9B9A9875B5;
defparam prom_inst_2.INIT_RAM_3F = 256'h9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9ABABBBB08EBEB;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[23:0],dout[31:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 8;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h3E3E3A3E423E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E;
defparam prom_inst_3.INIT_RAM_01 = 256'h46464A4A423E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E;
defparam prom_inst_3.INIT_RAM_02 = 256'h3E42423E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E;
defparam prom_inst_3.INIT_RAM_03 = 256'h46464A4A464A423E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E424242;
defparam prom_inst_3.INIT_RAM_04 = 256'h424646423E424242424242424242424242424242424242424242424242424242;
defparam prom_inst_3.INIT_RAM_05 = 256'h4A4A46464A4A464646423E424242424242424242424242424242423E3E424246;
defparam prom_inst_3.INIT_RAM_06 = 256'h42191D4246424246424242424242424242424242424242424242424242424242;
defparam prom_inst_3.INIT_RAM_07 = 256'h4A4A464A4A4A4A4A4A4A464242424242424242424242424242424642463A1525;
defparam prom_inst_3.INIT_RAM_08 = 256'h05120A254E463E3A464A42424242424242424242424242424242424242424242;
defparam prom_inst_3.INIT_RAM_09 = 256'h4A4A4A4A4A4A4A4A4A4A4A4242424242424242424242424642463A3E42111209;
defparam prom_inst_3.INIT_RAM_0A = 256'h090A0E1532250905213646424242424242424242424242424242424242424242;
defparam prom_inst_3.INIT_RAM_0B = 256'h4E4E4A4A4646464646464646424242464A46424242424242462E0D1919051212;
defparam prom_inst_3.INIT_RAM_0C = 256'h0501160E0505160E01092E4A4242424242424242424242424242424242424242;
defparam prom_inst_3.INIT_RAM_0D = 256'h4A4A4A423A363A3A3E42424242424A4E4E4A4A464242424636050E09050A0A0D;
defparam prom_inst_3.INIT_RAM_0E = 256'h12120E0E0E0A0E12161205364A42424242424242424242424242424242424242;
defparam prom_inst_3.INIT_RAM_0F = 256'h4E4A3E36363636363A3E42464A4E4E4E4E4E4E4E46424A3A0912120A0F13120D;
defparam prom_inst_3.INIT_RAM_10 = 256'h0E130F0E12130E0E1212012D4A42464646464646464646464646464646464646;
defparam prom_inst_3.INIT_RAM_11 = 256'h4E423636363A3A3636363A424E4E4E4E4E4E4E4E4A4E5225010E0E0E120E120F;
defparam prom_inst_3.INIT_RAM_12 = 256'h0E120F12120E0E0E05010D3A4642464646464646464646424246464242424646;
defparam prom_inst_3.INIT_RAM_13 = 256'h3E363636363A3A3636363636464E4E4E4E4E4E4A4E5B32051209120F12120A0E;
defparam prom_inst_3.INIT_RAM_14 = 256'h16130B0E12120E0911052152464A464646464646464646464646464646464646;
defparam prom_inst_3.INIT_RAM_15 = 256'h36363636363A36363636363636464E4E4A4A4E4E4F2E0109120E0A120E0F1215;
defparam prom_inst_3.INIT_RAM_16 = 256'h0A060A0A120F0E120A05093A57524E4A46464646464646464646464646464646;
defparam prom_inst_3.INIT_RAM_17 = 256'h3636363636363636363636323636424A46464A4A4A150A0D0912120E0E050E12;
defparam prom_inst_3.INIT_RAM_18 = 256'h0E0E16130E0E0E11090A092546574E4E4A4A4642464646464646464646464646;
defparam prom_inst_3.INIT_RAM_19 = 256'h3636363636363636363636363636363A4646462A08051212050A0F12160D0E0B;
defparam prom_inst_3.INIT_RAM_1A = 256'h13130E120A0A0E0D1205090501365353524A4646464646464646464646464646;
defparam prom_inst_3.INIT_RAM_1B = 256'h363636363636363636363636363636363E4642040905090E13130E170E0E1212;
defparam prom_inst_3.INIT_RAM_1C = 256'h0E0A0E0D0E12120F0A06160E011953534F4E4E534E4646464646464646464646;
defparam prom_inst_3.INIT_RAM_1D = 256'h36363636363636363636363636363636363A422905050109120E0E0A0E160E12;
defparam prom_inst_3.INIT_RAM_1E = 256'h12050E0E120E0E060E1312091D4A534F4E4F534F4E4A46464646464646464646;
defparam prom_inst_3.INIT_RAM_1F = 256'h3636363636363636363636363636363636363A521D011105090E120A0E120A0E;
defparam prom_inst_3.INIT_RAM_20 = 256'h0A0E120A130B0E160D0E090036574A4E4E4A4E4A4A4A4A4A4A46464646464646;
defparam prom_inst_3.INIT_RAM_21 = 256'h3636363636363636363636363636363636363A320409090905090E0A0E0E120F;
defparam prom_inst_3.INIT_RAM_22 = 256'h12120F0A0E1216120509090D04314A4A4A4A4A464646464A4A4A4A4A4A46464A;
defparam prom_inst_3.INIT_RAM_23 = 256'h3636363636363636363636363636363636363A361901050909110D050E12120E;
defparam prom_inst_3.INIT_RAM_24 = 256'h090A12120909110909090909051D4E4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4F;
defparam prom_inst_3.INIT_RAM_25 = 256'h36363A363636363636363636363636363636363611010D0E0D0E120E0E0E0F0E;
defparam prom_inst_3.INIT_RAM_26 = 256'h090911110A0E010512160E010D424A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4E5353;
defparam prom_inst_3.INIT_RAM_27 = 256'h36363A363636363636363636363636363636362A000505050505090E0A0A0E09;
defparam prom_inst_3.INIT_RAM_28 = 256'h0E0E1212160E09090E0A010901194F4A4A4A4A4A4A4A4A4A4A4A4A4F53535353;
defparam prom_inst_3.INIT_RAM_29 = 256'h36363636363636363636363636363636363636320D05091609090E120D12120E;
defparam prom_inst_3.INIT_RAM_2A = 256'h0E1612050901091205050501083A4F4A4A4A4A4A4A4A4A4A4A4A4F5353535353;
defparam prom_inst_3.INIT_RAM_2B = 256'h363636363636363636363636363636363636363E1D00090A050E0E050D05090E;
defparam prom_inst_3.INIT_RAM_2C = 256'h090D050D090D120E090D0D0036534A4A4A4A4A4A4A4A4A4E4F53535353535353;
defparam prom_inst_3.INIT_RAM_2D = 256'h3636363636363636363636363636363636363636360D050505090905090E0505;
defparam prom_inst_3.INIT_RAM_2E = 256'h0905091109090909050100114A4F4A4A4A4A4A4A4A4F4F535353535353535353;
defparam prom_inst_3.INIT_RAM_2F = 256'h36363636363636363636363636363636363636363E1D0004050D0901090E0509;
defparam prom_inst_3.INIT_RAM_30 = 256'h0D0505050905090909212146574E4F4F4F4F4F4F4F4B4F5353534F4F4F535353;
defparam prom_inst_3.INIT_RAM_31 = 256'h3636363636363636363636363636363636363636363E21110109010005090805;
defparam prom_inst_3.INIT_RAM_32 = 256'h050405090D05080109575B534B4B4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F;
defparam prom_inst_3.INIT_RAM_33 = 256'h363636363636363636363636363636363636363636363E361508363A19142009;
defparam prom_inst_3.INIT_RAM_34 = 256'h0C1C0D05001D320D3A534F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F;
defparam prom_inst_3.INIT_RAM_35 = 256'h36363636363636363636363636363636363636363636363A36324A5B4E253D1C;
defparam prom_inst_3.INIT_RAM_36 = 256'h28311C0D194A5353534F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F;
defparam prom_inst_3.INIT_RAM_37 = 256'h3636363636363636363636363636363636363636363636363636363E4F294535;
defparam prom_inst_3.INIT_RAM_38 = 256'h353514315B534F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F53534F4F;
defparam prom_inst_3.INIT_RAM_39 = 256'h363636363636363636363636363636363636363636363636363636363A295145;
defparam prom_inst_3.INIT_RAM_3A = 256'h41391C39574F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F534F4F4F4F46424236;
defparam prom_inst_3.INIT_RAM_3B = 256'h36363636363636363636363636363636363636363636363636363A3632255A49;
defparam prom_inst_3.INIT_RAM_3C = 256'h412D312842534F4F4F534F4F4F4F4F4F4F4F4F4F4F534F463A3A3A3A36362E26;
defparam prom_inst_3.INIT_RAM_3D = 256'h3636363636363636363636363636363636363636363636363636363636215555;
defparam prom_inst_3.INIT_RAM_3E = 256'h4124352842574F5757465B5357534F4F4F4F53534B463E3636363636362E262A;
defparam prom_inst_3.INIT_RAM_3F = 256'h36363636363636363636363636363636363636363636363636363A3636255955;

endmodule //Gowin_pROM
